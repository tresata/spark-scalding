name|color|quantity
apple|red|5
grape||50
pear|green|3
